//*****************************************************************
//*	描    述:	待测信号输入缓存
//*	开始时间:	2015-03-14
//*	完成时间:	2015-03-14
//*	修改时间:	2015-03-15
//*	版    本:	V1.0
//*	作    者:	凌智电子
//*	说    明:	使待测信号与系统时钟同步
//*	备    注:	
//*****************************************************************

module in_buf (
	input  clk,			// 驱动时钟
	input  in_a,		// 待测输入信号 a
	input  in_b,		// 待测输入信号 b

	output q_a,			// 同步后输出信号 a
	output q_b			// 同步后输出信号 b
);
// 信号a缓存寄存器
reg                        ina_r = 1'b0;
// 信号b缓存寄存器
reg                        inb_r = 1'b0;


//*****************************************************************
//* 待测信号输入一级缓存, 使其与系统时钟同步
//*****************************************************************
always @(posedge clk) 
begin
  ina_r <= in_a;
  inb_r <= in_b;
end

assign q_a = ina_r;
assign q_b = inb_r;

endmodule 

//*****************************************************************
//*                    END OF FILE 
//*****************************************************************