//*****************************************************************
//*	描    述:	待测信号异或
//*	开始时间:	2015-03-14
//*	完成时间:	2015-03-14
//*	修改时间:	2015-03-15
//*	版    本:	V1.0
//*	作    者:	凌智电子
//*	说    明:	使待测信号异或输出, 其它控制信号需一级缓存, 保证输
//*			出同步. 
//*	备    注:	
//*****************************************************************

module buf_or (
	input  clk,			// 驱动时钟
	input  rst_n,		// 复位信号
	input  ina,			// 待测信号 a 输入
	input  inb,			// 待测信号 b 输入
	input  o_en,		// 闸门控制信号输入
	
	output ina_out,	// 待测信号 a 输出
	output inb_out,	// 待测信号 b 输出
	output cnt_en,		// 闸门控制信号输出
	output q				// 异或输出
);

reg  [1:0]	cnt_en_r = 2'b00;
reg         q_or = 1'b0;
reg  [2:0]  ina_r = 3'b000;
reg  [2:0]  inb_r = 3'b000;


//*****************************************************************
//* 待测信号异或
//*****************************************************************
always @(posedge clk) 
begin
	q_or <= ina ^ inb;
end

assign q = q_or;

//*****************************************************************
//* 闸门控制信号缓存
//*****************************************************************
always @(posedge clk) 
begin
	cnt_en_r <= {cnt_en_r[0], o_en};
end

assign cnt_en = cnt_en_r[0];

//*****************************************************************
//* 待测信号 a 缓存
//*****************************************************************
always @(posedge clk) 
begin
	ina_r <= {ina_r[1:0], ina};
end

assign ina_out = ina_r[0];

//*****************************************************************
//* 待测信号 b 缓存
//*****************************************************************
always @(posedge clk) 
begin
	inb_r <= {inb_r[1:0], inb};
end

assign inb_out = inb_r[0];

endmodule 

//*****************************************************************
//*                    END OF FILE 
//*****************************************************************